library ieee;
use ieee.std_logic_1164.all;

entity reg is
    generic (width: integer := 8);
    port (
        clk: in std_logic;
        resetn: in std_logic;
        loadEnable: in std_logic;
        dataIn: in std_logic_vector(width-1 downto 0);
        dataOut: out std_logic_vector(width-1 downto 0)
    );
end entity reg;

ARCHITECTURE behaviora OF reg IS 
BEGIN

  PROCESS ( clk , resetn ) 
  BEGIN
    
    IF resetn = '0' THEN
    	dataOut <= (OTHERS => '0');
    ELSIF rising_edge(clk)THEN --(rising_edge(clk) AND loadEnable='1')
	IF loadEnable='1' THEN
		dataOut <= dataIn ; 
	END IF;
    END IF ;

  END PROCESS ; 
END behaviora;